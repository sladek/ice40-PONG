/**************************************
* Module: character_memory
* Date:2018-04-29  
* Author: sladekm     
*
* Description: 
***************************************/
module  character_memory(
    input   [7:0]  address,
    output  reg [7:0]   data
);


always @*
  begin
     case(address)
// 0 - '0'
       8'd0 : data =  8'b00011110;
       8'd1 : data =  8'b00100001;
       8'd2 : data =  8'b00100001;
       8'd3 : data =  8'b00100001;
       8'd4 : data =  8'b00100001;
       8'd5 : data =  8'b00100001;
       8'd6 : data =  8'b00100001;
       8'd7 : data =  8'b00011110;
// 1 - '1'
       8'd8 : data =  8'b00000010;
       8'd9 : data =  8'b00000010;
       8'd10 : data = 8'b00001110;
       8'd11 : data = 8'b00000010;
       8'd12 : data = 8'b00000010;
       8'd13 : data = 8'b00000010;
       8'd14 : data = 8'b00000010;
       8'd15 : data = 8'b00000010;
// 2 - '2'
       8'd16 : data = 8'b00011110;
       8'd17 : data = 8'b00000001;
       8'd18 : data = 8'b00000001;
       8'd19 : data = 8'b00011110;
       8'd20 : data = 8'b00100000;
       8'd21 : data = 8'b00100000;
       8'd22 : data = 8'b00100000;
       8'd23 : data = 8'b00011110;
// 3 - '3'
       8'd24 : data = 8'b00011110;
       8'd25 : data = 8'b00000001;
       8'd26 : data = 8'b00000001;
       8'd27 : data = 8'b00000110;
       8'd28 : data = 8'b00000001;
       8'd29 : data = 8'b00000001;
       8'd30 : data = 8'b00000001;
       8'd31 : data = 8'b00011110;
// 4 - '4'
       8'd32 : data = 8'b00100000;
       8'd33 : data = 8'b00100010;
       8'd34 : data = 8'b00100010;
       8'd35 : data = 8'b00011111;
       8'd36 : data = 8'b00000010;
       8'd37 : data = 8'b00000010;
       8'd38 : data = 8'b00000010;
       8'd39 : data = 8'b00000010;
// 5 - '5'
       8'd40 : data = 8'b00011111;
       8'd41 : data = 8'b00100000;
       8'd42 : data = 8'b00100000;
       8'd43 : data = 8'b00011110;
       8'd44 : data = 8'b00000001;
       8'd45 : data = 8'b00000001;
       8'd46 : data = 8'b00000001;
       8'd47 : data = 8'b00111110;
// 6 - '6'
       8'd48 : data = 8'b00011110;
       8'd49 : data = 8'b00100000;
       8'd50 : data = 8'b00100000;
       8'd51 : data = 8'b00111110;
       8'd52 : data = 8'b00100001;
       8'd53 : data = 8'b00100001;
       8'd54 : data = 8'b00100001;
       8'd55 : data = 8'b00011110;
// 7 - '7'
       8'd56 : data = 8'b00111110;
       8'd57 : data = 8'b00000001;
       8'd58 : data = 8'b00000001;
       8'd59 : data = 8'b00000110;
       8'd60 : data = 8'b00001000;
       8'd61 : data = 8'b00001000;
       8'd62 : data = 8'b00001000;
       8'd63 : data = 8'b00001000;
// 8 - '8'
       8'd64 : data = 8'b00011110;
       8'd65 : data = 8'b00100001;
       8'd66 : data = 8'b00100001;
       8'd67 : data = 8'b00011110;
       8'd68 : data = 8'b00100001;
       8'd69 : data = 8'b00100001;
       8'd70 : data = 8'b00100001;
       8'd71 : data = 8'b00011110;
// 9 - '9'
       8'd72 : data = 8'b00011110;
       8'd73 : data = 8'b00100001;
       8'd74 : data = 8'b00100001;
       8'd75 : data = 8'b00011110;
       8'd76 : data = 8'b00000001;
       8'd77 : data = 8'b00000001;
       8'd78 : data = 8'b00000001;
       8'd79 : data = 8'b00011110;
// 10 - ' '
       8'd80 : data = 8'b00000000;
       8'd81 : data = 8'b00000000;
       8'd82 : data = 8'b00000000;
       8'd83 : data = 8'b00000000;
       8'd84 : data = 8'b00000000;
       8'd85 : data = 8'b00000000;
       8'd86 : data = 8'b00000000;
       8'd87 : data = 8'b00000000;
// 11 - '-'  
       8'd88 : data = 8'b00000000;
       8'd89 : data = 8'b00000000;
       8'd90 : data = 8'b00000000;
       8'd91 : data = 8'b00111110;
       8'd92 : data = 8'b00000000;
       8'd93 : data = 8'b00000000;
       8'd94 : data = 8'b00000000;
       8'd95 : data = 8'b00000000;
// 12 - 's'  
       8'd96 : data =  8'b00000000;
       8'd97 : data =  8'b00000000;
       8'd98 : data =  8'b00000000;
       8'd99 : data =  8'b00000110;
       8'd100 : data = 8'b00001000;
       8'd101 : data = 8'b00000100;
       8'd102 : data = 8'b00000010;
       8'd103 : data = 8'b00001100;
// 13 - 'L'  
       8'd104 : data = 8'b00000000;
       8'd105 : data = 8'b00000000;
       8'd106 : data = 8'b00000000;
       8'd107 : data = 8'b00001000;
       8'd108 : data = 8'b00001000;
       8'd109 : data = 8'b00001000;
       8'd110 : data = 8'b00001000;
       8'd111 : data = 8'b00001110;
// 14 - "live" symbol  
       8'd112 : data = 8'b00000000;
       8'd113 : data = 8'b01101100;
       8'd114 : data = 8'b11111110;
       8'd115 : data = 8'b01111100;
       8'd116 : data = 8'b00111000;
       8'd117 : data = 8'b00010000;
       8'd118 : data = 8'b00000000;
       8'd119 : data = 8'b00000000;

// 15 - 'G'  
       8'd120 : data = 8'b00111110;
       8'd121 : data = 8'b01000001;
       8'd122 : data = 8'b01000000;
       8'd123 : data = 8'b01000000;
       8'd124 : data = 8'b01001111;
       8'd125 : data = 8'b01000001;
       8'd126 : data = 8'b01000001;
       8'd127 : data = 8'b00111110;

// 16 - 'A'  
       8'd128 : data = 8'b00001000;
       8'd129 : data = 8'b00010100;
       8'd130 : data = 8'b00100010;
       8'd131 : data = 8'b01000001;
       8'd132 : data = 8'b01111111;
       8'd133 : data = 8'b01000001;
       8'd134 : data = 8'b01000001;
       8'd135 : data = 8'b01000001;

// 17 - 'M'  
       8'd136 : data = 8'b01000001;
       8'd137 : data = 8'b01100011;
       8'd138 : data = 8'b01010101;
       8'd139 : data = 8'b01001001;
       8'd140 : data = 8'b01000001;
       8'd141 : data = 8'b01000001;
       8'd142 : data = 8'b01000001;
       8'd143 : data = 8'b01000001;

// 18 - 'E'  
       8'd144 : data = 8'b01111111;
       8'd145 : data = 8'b01000000;
       8'd146 : data = 8'b01000000;
       8'd147 : data = 8'b01111000;
       8'd148 : data = 8'b01000000;
       8'd149 : data = 8'b01000000;
       8'd150 : data = 8'b01000000;
       8'd151 : data = 8'b01111111;

// 19 - 'O'  
       8'd152 : data = 8'b00111110;
       8'd153 : data = 8'b01000001;
       8'd154 : data = 8'b01000001;
       8'd155 : data = 8'b01000001;
       8'd156 : data = 8'b01000001;
       8'd157 : data = 8'b01000001;
       8'd158 : data = 8'b01000001;
       8'd159 : data = 8'b00111110;

// 20 - 'V'  
       8'd160 : data = 8'b01000001;
       8'd161 : data = 8'b01000001;
       8'd162 : data = 8'b01000001;
       8'd163 : data = 8'b01000001;
       8'd164 : data = 8'b01000001;
       8'd165 : data = 8'b00100001;
       8'd166 : data = 8'b00010010;
       8'd167 : data = 8'b00001100;

// 21 - 'R'  
       8'd168 : data = 8'b01111110;
       8'd169 : data = 8'b01000001;
       8'd170 : data = 8'b01000001;
       8'd171 : data = 8'b01111110;
       8'd172 : data = 8'b01001000;
       8'd173 : data = 8'b01000100;
       8'd174 : data = 8'b01000010;
       8'd175 : data = 8'b01000001;

       
// Default
       default : data = 8'b00000000;
    endcase
end 

endmodule

